timescale '1ns/1ns


module ();

endmodule
always @(posedge clk or negedge rstn) begin
    
end